class transaction;
  randc bit a;
  randc bit b;
  randc bit cin;
  bit sum;
  bit carry;
endclass
