interface segment_if;
  
  logic [3:0] bcd;
  logic [7:0] segment;
  
endinterface
