class transaction;
  randc bit a;
  randc bit b;
  
  bit difference;
  bit borrow;
endclass
