interface hs_if;
  logic a;
  logic b;
  logic difference;
  logic borrow;
endinterface
