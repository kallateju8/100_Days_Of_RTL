interface transmission_if;
  logic a;
  logic control;
  logic y;
endinterface
