interface demux_if;
  logic d;
  logic [1:0]sel;
  logic [3:0]y;
endinterface
