class transaction;
  randc bit a;
  randc bit control;
  logic y;
endclass
