class transaction;
  rand bit d;
  rand bit [1:0]sel;
  bit [3:0]y;
endclass
